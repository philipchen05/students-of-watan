Blue
0 0 0 0 0 g c 1 1 23 1
0 0 0 0 0 g c 2 1 19 1
0 0 0 0 0 g c 6 1 15 1
0 0 0 0 0 g c 8 1 11 1
4 3 4 10 0 11 4 4 2 5 0 8 1 3 2 11 5 7 3 10 3 12 2 9 3 9 0 5 1 8 1 2 0 6 1 6 2 4
-1

Blue
999 1999 2999 4000 4999 g 44 39 31 22 c 0 3 33 3 26 3 14 1
0 0 0 0 0 g c 9 1 37 1
1 0 0 0 0 g c 11 1 48 1
0 1 0 0 0 g c 24 1 45 1
4 3 4 10 0 11 4 4 2 5 0 8 1 3 2 11 5 7 3 10 3 12 2 9 3 9 0 5 1 8 1 2 0 6 1 6 2 4
8
